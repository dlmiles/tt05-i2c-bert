//
// SPDX-FileCopyrightText: Copyright 2023 Darryl Miles
// SPDX-License-Identifier: Apache2.0
//

//
//
//


`ifndef SYNTHESIS_OPENLANE
`ifndef UNIT_DELAY

//`define UNIT_DELAY

`endif 	// UNIT_DELAY
`endif	// SYNTHESIS_OPENLANE
